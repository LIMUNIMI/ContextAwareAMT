BZh91AY&SYIm*W_�|x���������a7�>
>}1�(@H`
 
)J`                                �
U >       �| �                  �                  �   �$�$@D��!@:�D�   тU_ 4P��*ADTD�  �)� �   | �*B
��� 	Ѕ	 �T�  �    ����鈄
DB �{i��p �J�  @ �   � ,�I  "$;2���P�   �   �J�@��B��P
���@  � �   8TEJ�� �� �*�R�R���$=  S�  �`�^$Q'�  � T�@   p   $�($H�  g ( "U �"��$@"�*�#�        j���)T����~�  �  U6ު�U2adi�@��4ш4h���J��=�z��4�@�����bOU*���h      �T����M4�*6�=�yOMO�<���T��ҁU?T�������UR��@      ��}����>�}�w��HE^i?����H��QIO��*���_��ľ�/�_?7��^K�y/%���x�x�x�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x�����������9�9�9��<s�<s�<s�<s���y/%众����^K�y/%�9�s�<s�<s�<s�=�x�x�x�x�����������9�9�9��y��w��;rctr���[t�c]#���K�c9�|]lDGN" ��Y��&X�����g9c��M���
(�8�QN�b���1vQEӱH�^���{Μ���s�<s�<s��x�x�x�{���������{�9�9�9�9�s�<s�众��^|�K�y/%众����9�9�9��<s�<s�<���^z��7��^K�y/%��x�x�x�x�����������9�9���>9�ϋ�^������^K�y/%众�����������9�9�9��<s�<s�<s�<s��x�x�x�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x�����������9�9�9��<s�<s�<s�<s��x�x�x�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x����^K�y/%��众��^K�<s��x�x�x�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x�����������9�9�9��<s�<s�<s�<s��x�x�x�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x�����������/%众��^|�K�y/%众�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x�����������9�9�9��<s�<s�<s�<s��x�x�x�{���������{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x�����������9�9�9��<s�<^K�y/%��众��^K�y/{�9�9�9�9�s�<s�<s�<s�=�x�x�x�x���^K�y/%���"��|�������L3BE^ ������/@��م��{d�������x=���i�_�鴶M�kd-&-��j64E��ccDX��6%mVV��-��j1�V5V+&-��Z-�j4E��ccDZ*"�P*��X�Z��(ڍ�cj6�6�cb����E��-h��EDkS&ȶkj6�j2�U�m���6ƍ�E��Q�F�V-E��h�h�E��1Eb�(�Q�(�1�Q�c�1�c�1�c�1��������������,h�M�ƭb��m�TkJ��6�����h�Z-�F��QQQQQQQQQ�cE�,h�cFō,h�՚�ؓeM�d0��klk�cX�k�F�h�Z-�F�������Ŋ��
��E�&�l��VjM���j6���6���b�X�Z-���h�%��l%m+T���hڋQ�b��b��6�E��h�m	�ʖ�[)�V�[R��kk*6���X�Z1�h�Z-�E����4E4XѢƍ
&�i�H6��&�+�+ƣu������us���y�o��z�w�=���<��G����o��z=��G�Ę�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�|��k�Ϛֱ�I�cĘ�1��5�c�ֵ�c��kX��1�1�c�ֵ�~kZ�1��kX�Ϛֱ�|��kĘ�1�I�c��Z�1��kZ�>|ֵ�1�cc�1��kX�浭c�ֵ�<���y6�N������:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t���:GH�#�t����:GH�#�t���":GH�#�t���:GH��#�t���:GH�"#�t�1�8��z�z�^�_����/瞏C���y�z�~?�{��5�w��7��zR�x���~�-�vM��v���SƓ�^5Ge�[ض*ŬZ5F��Ej-���-cm�\��F�Ɠ�Sb�V�/�Fʿvh�&�lma���lW�Q�Cj5�m�b�ZţTml�b;+�lVҶV�-��;*�6��&Ľ1ڍ��l�-��Gev*�����.�vN�66��6�حElj-�Z��lj*���EU�ca�I���V���mFʻ�M�e66���Si6+�TvP��VʶV���Cƥv��b���+�Kc�Fʹ\U��E���6���el�b�Q��v�����[I�;$��W��kb����5kj-�F�ګd���Q�v��Tm�lj�(ڋm�]�l�)��-�ʛI�]�=2��i^2���]��6�ԭ��l��b�����lmQ�*�l-��6%��Q�l�evK�ڍ��VжU�i<d�ci]�`�[�[F��%��*�;�V����6���ح����V������ݟ?	~��?��ﾾ�������������         lxG��                                         ��????                                                                w  =�                                                    ���                                                                                                                      �`                                                                                        �������U����|�E_�������m�i�Q���wwwwwwwwr���������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_''�������_��W�B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!o���E__T%i�m�W*�u�  2L� �2  $� �2  $�d �L� �I� L� I&@ I2  $�  2I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$��I$�$I$�I2H�I$�d�$�I$ȒI$�d�$�I$ȒI$�dI$�I2$�I$�I$�L�$�I&D�I$�&I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�RI$�I#̻���fg񙙙�m���H�I$�I�0�  KZI$I"I$���m�   5�I$�$I$�s0  �`��$�I$�D��  ��Z�I$�I$�[�`��m�  -t�$�I$�.a�m� m��֒IH�I/nn�    k��IH�I>�0`� l>�H�I$�Il6� ��KZI$I"I$�� ��l ��I$I"I$���`   6���I$�I$�9���   u�ZI$�I$�K{   m�� Z�I$�I"\� �  ���H�D�I{v��`  ]$�H�D�I�0   �`��$�I$�D��   m�:��$�I$�I%�� �m�  -t�$�I$�&��  �KZI$I"I$�s�    t�I"II%�f �����$�I$�D�f  6� �n�kI$�I$�I��m��   ��$�I$�$�  � �֒IH�I-ݘ   m���$�$�$�]�`m��� �]"I$�I$K�`� 6� �ִ�I$�I$�f�    ��$�I$�$���  ��kI$�$I$���  �m��$�D�$�O���   �]"I$�I$K���� ׭i$�I$�I>��   6�k��I$�I$�6`  �`��$�$�$�[�0 m��  k��IH�I.�6�   ��u�I$�I$K�a��   u�ZI$�I$�O�0  6�m�-t�$�I$�&� m� ��$�$�$�[�1��l   k��IH�I.�0  m�>�H�I$�Is   ���ִ�I$�I$�� m��  ��$�I$�D��m�  m�zZ�I"II%�Ͱ    k��IH�I>�  m����t�$�I$�'0  m���z֒I$�I$�����l   �D�I$�H��  6� KZI$I"I$��    m׭i$�$�$��`l m� >�H�I$�Is l m�׭i$�I$�I-��    ]"I$�I$K� 6�  6޵�$�$�$�^݀  6�m��I$�$�$�|� 6�  ��I$�I"Nm� 6�  :��$�I$�I%��   ���I$�I"\��  � =-i$�$�$��� �m� �I$�$�$��cm�   ���$�I$�$��   ׭i$�I$�I-�  ��lk�I$�I$�s  6�  zZ�I"II%��6�m�  t�I"II'��  m�>�H�I$�Is   ���ִ�I$�I$�� m��  ��$�I$�D��m�  m�zZ�I"II%�Ͱ    k��IH�I>�  m����t�$�I$�'0  m���z֒I$�I$�����l   �D�I$�H��  6� KZI$I"I$��    m׭i$�$�$��`l m� >�H�I$�Is l m�׭i$�I$�I-��    ]"I$�I$K� 6�  6޵�$�$�$�^݀  6�m��I$�$�$�|���m�  }��$�I$�$�ݱ�m�  u�ZI$�I$�K{  ��]u�I$�I$K��  l ����D�$�K۱���l ��I$I"I$���`   6���I$�I$�9�n�   �kI$�I$�Iw�}_H�$�����Y�+Y[m�-2��,+R��J�,��YxV��j�%��ҥ��ж�Q���[,�V�m��X�2�V���JZ$e�XV����jYe���E��-8K,	e�Kem�R��/,��Z��lF��X��ңmBӄ��,��ֵ��Rв�2�V����ae��Z��ڍ-���e�Km����X��R����R�#/,�µ-���R�,�%��j-��i�Y`K-*[+m���Yye�
�V�b4����V��j�%�Ye�6���Җ��X��R�m����-�X��-��ile��(�[mE��2Ō�����Җ�ye��mm�Z�Ye�,�+Qm�N�YiR�[l����,�V����%������P��,��,���m���,�Ō���m��XFYl��֩m��Kc,�Y@�R�j-l���m-��<,*R5^Z�,����-c
��(QB��"2�兖[/-(�+i���!Bլo,����KQ%![K[b�-m�R�,�������<�w������}g�?�6駍/���O��R��X���V}�Oz��붬i�M7 �x�n��]�O.�>�u�ޯ�w����HcH1t�,f��m�ҷJ;X[2����;�����d�+׿]����O|�Nrkλ.�ޖm�v=+�{��36���W�$�k3]�ґ���Y���qnJ�$�]�y���߻�I�O����OD7Gk��a%��ْ]H�[��뵵3o�{f��Un������m�[���֙����]v�p_}��I��6�E��H�"khyC���^�����}���+z����u/���ye��u6�s��@��:�Z�;�������=��l=ml��;�{8=��,�iq��d�­�,M9�i�mpw���}�v�w�W��D�������a����e����ΚG5�q�5�1o5ǝ��ow�o2D�ɝ���vYNՙ&fL�nono�rDl�}�q��j}������Gjk#����r�>�i�D�97}���r�n^��i�Y�hm���Sf����N`��˭�j�fC<�t�]lQ�K]��؄�\L�t˙�&����a���\j��ɝ�H.��[4�S;��d�R�-�,�%�y����6s��Me]n�8�4�w1[��H����ǹ�ۻ�[��k�s��}G#�m�O����U��5בI:�wj8�:<�s�|"
n}�R���]a������Z�}�w���ܕ�M�ؙ3#�mo_%�ʭ���E��6��kzf�u �����N,��fϳRN��󱾝5ζ�Zyn*��]�+���w��e�췸��)Z�ɧ����4wwDrjIɍvI6�w��c��k��D��rL�oQ���'	��s��M�93��>m�|�����Ue�|�I�G�['RDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDHI���g����>��5�]��\�3r1V�����6v����um;�=V�m6�.M8��Iw��w�VA9�Oo�)w���"�f�-=C�1�Y;�v�/$�98^�~|b�����<g��Ԟn��)�as��.�۩���d�)��amk6�����z�w~����w���f9׾�'_=��co���H���4�#�T�OSX�F�/�^<;{��L�}�s�s����w�[�;�$����_�'���n^&��ҙ�uXV��,a��2.�ɳ`YV��I�nL�ʺ�nR��fe�3��GXQ�n�n�k�� 0bd�e���8@бt.a�s��vaSV9�l�q4tD�nFz�3�o��1�N�e��]�R�oWy�>�o���a��)S��3�����}���l�ck������gޏ}���>�=]�;y����z@��׶����opܺ���5�M��ZjfH��)Slh���@�ܖ]��S.��f�[��[�ޔ���xɮ�o���L�LZd�۵q�����oL�];r�S��տ�$��/#�$��i��'b�o!_�wa�O~�|�U���h�*����K���6��LE����λ�K��m.v����ɧv�5�qL��yd��7��Kh��������A���1�A� �ac0�A�� �a0�1�A� �ac0�A�� �rs������3��55��x�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0���+�_�+�/�U��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU^y�y�y������8�����	G����Q�'8�;���K�]s�s�"��$��4��-�]��k��~y$b�C�Q���/�\_��gǛgt��|��<���5�M����.���&�f�We�B${���~�{�s����d�_�q��T�|�s�}��'@ygd�?�I9�NNr~�:��Y��N�����w�s���I��M�񪥣��'}�)��I/�N���\��>u����&=��=�w/Vۿ���g�ً�$��)��������.m���q �*�ަy��y��_�Y�z_��V\���Cw�����O�=�)�����Y�o���hҍ�Ż&���{�fdqe�_�I9�tc�������~����}P��3�ϯ��n������y���{g�����3$m%��W�K����<mmx=$5��k�P��.&X���#��6���)��I�`�u���b�S,]A�(�J�mL�1�	0�
i�f�%����l9ٔՖ�sq�a�o+�Ώ,�qv���s2`����R[�����l����pBi�o�K�d�wO�wS,���N6��$��W�R~��i�r޹ĝ�9=ts�A	�rtN':'�yy:'+;!���ٔ�I�C���m�y��!�brK<h�oK9Z���s��8��s)���v�u�+?u�Ǎnĺ�H�4�k��0��sYvj���߻�'��AS�����Jtc�\Oo~A���C�'�<�2BBHHH�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"����)�Z����ln������U��l�n�g����}f'���V���NruN���i�tu��߻�*���Z�.�[���~;;�����}e%��?zO<�y��mWO�ݧR�׫��+�Yt�[E�y�-i>�:������¯��������q;u�O��Zjn,kÙȶ5��&^[2ez�^}�dz_-�d�s�����km���M��fk�k����=��4t�y������.���[��}�t���_��oК�LW�u�ٷ[M0M�6���a{����oGW��y���3�^{|���s��+�I��ӯ��>b��y�?>B�=��S��{n�Ǿ�_��q�cOjK#�%�QwsN�g���m��=~E�:����9�����韑_g7w̳Λ=�3|z{/�᭺h-��Wit��6��f�M��Yו�{������C�2vD�7z�-{믙:$��~~�������r�KY�%%�P�䤞O��w%'��O��c�QD�_|�>3�Mr�x��MF��v,D�;5w�ZY�ǽ����H����%�N������jś��w���}u��ɤ6��F�e+�p��X�Ch02h�kv�\�bMɸh.�$6n&.�1̱ԃ��b�+M�6L�8��!�0R��Mv�	N h;9nU�̺[,�X��FfL#9.��� ���K�fnF*�@5�l���9��S��ۉ���?�e>�ZϞv�ꐛ�x�R~�:�����n�3�׽Lȍ�<xץޑٵ�֥�o>��w�[k��dW5�7���Y���?w[�#��ưe"O�f6��oR���G��΍�7���ļ����!s��ˁ��Sbg:2d�uѬ�f��ߵ�������2V�"M�M���z)�����Z�nrI/�^I%��-?��jg�[�~^g����g�v�5��O�I%��}���~Y~~&���������w��\W�s�|޹�¾��H�d�����XM���7�����2wƷb]pP&�it�g:a[���k����ST�3��:�����|�"�&f��53[����؏rI�kY;,|������교iؓ�nF�M�y�_W�z3�[�7�xY���3�ޟo��&�ܑ��ˋ���y��/�#hh[��k�����n���������9|rxtI�N��G��z�;χ~O��R�{�~�trC�vt,kw�}��u�7#̞o�����_|�X��g��I/�S�z}��e�k��=f�F����q-8�ɷ=~nu���4��o�r�������y��=9�[[E��5���.�Y]�p5���t���|w��\U������n.nkZ��+���*����{�~�տ��y�diG��g�3�z�\�ȷ�>�z�1Ď7]ޱ��,7���{ϸ��1m�X����[��V��ߛ����3���b������o�?����a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�������VɴUm[Kb5V5�F-���F�-��ر�6,h��#bƈ�Z׉U��mF���m������X�جb�Q���TE��-��Sa6M�mVcj6�lmEcclm��l�E��hѢ�h�kw-�[T���i-�m4��liF�Y�i�ж��mKd���آ�Tأ4�Դ�"[*�	�"�Ƭ��բ�h�Z-(��h��QE��1Eb�1�c�1��1�c�1�c�"""1cE�4R��-�F��F�,TTT�H��،h���ƍ%�(��✥r�8�:�������<�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������P^B�z����k5�kSS���$��0s��|���%��9��;v�w������_����� �v��$��s��n��Z]�Iy�q��s�����s����9�Z���{��� �۝޺KޒX�/0]�s�zO�Kv��g9פ�u�1�v���s�]"I1�v���;�%��7m�y���9����i�9���nq-"I��9��v��%��t������;k�>I<�8��s�%�zIw��opݹ�뤽�%�r�۷9פ�$�m�y��s�zIw]#�n����=u�$��n���s��[Z�v���s��Z�֟c����v��$��s��n��Z]�Iy�q��s�����s����9�Z���{��� �۝޺KޒX�/0]�s�zO�Kv��g9פ�u�1�v���s�]"I1�v���;�%��7m�y���9����i�9���nq-"I��9��v��%����＂آ/nM�m��gJ�uf���L��]s6�q�&�``�ٸ��9U��@��v��&�9BMJ����$1 ó��15&��RgB�ɐÒ��"���t�5����.���ֻE������v?�_�ˉm�u���jF����Q�3���t��}�Kٶl��E�[�y��s;=Zj9
f�L�x���x\��o��6����}��1N��v�����]��J�_���S�IHˀ�@[�ՙv*��@5�6JgS��</���߿��ɻ��<�ٻ�i��;~)2�t~�+99���t�wKG_��I%�ˑnj��&9��������=��}1��c����v���gO�������,^j|����|4/4�I�YR��{+�I<��bIJ~��xs���L���:�!r�^2�mŸ�ؙΌ�0]w�t)e��G��ֲLs~Sﱫ�Ǧ�^�Ʈ�}��t\����}�'׉��y~��׫VzC��iF���i$��D��-�����*��]��I�2^#�i��w��bާÇ�u��s�_���=���S������QX�9מ\N�n��:�ƶ�fచ�.�l-�6k.��-n�y�첼���tw���:���K�8��^���y�s�{z���].m�=w��,��o��y^V��oX��}�C�ǟG�V,v��G�^��V�o"�L[k[�����w���/I;9�1�Os|�����O�e���x���S����gs�4-�Ե�h����@[HD��4�t���M�g��7�R���I2Mk��=�b�=������k�Ӎ{����fG��o��;�rxڋ��'�Eg$�nutU��۞�雙��^�C�f C��{z��a/E������戮s���;�TE��946ٗl�)t.Y�s�&L��]r\�ܛ���q��u�3�&6(����Sfbmr�75+���"�պ+�MHk�I��fd�Ò��m�Mcm1�ٵ�ٮ�ͦ���Q������9�f��޴�N�k\�ҧg��ܾ���N����c������[3%5�]�)�M{WzS'��K5w�ʛ�-�������'G>9O:��9N~9���F���i���G.e\_}��t����\���N�zS�����u����y���!�]�\��[���s�xJ��Iw|�Bv��q�~�ޣ�B'~9;�����ۯߞI�O�'�uqq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�qq�rq����������=9��ĥ��e��觢w:LOI�{����r��9{�qȬۑ?��c�t]%big\\k���_q���OBt_*=s�����
c����۴�wzC�M����"��.�˱UM��������$����Ϸgf�?�vt{z�����~������[��2^��Ӭk8��3$�m��C���Q����_ׂ7�L֢�̓�K����Sz�&'��[�}P�=9�m7+�Pq����d��e�55������jlL�<ɂ�U\��������������~��̓Y�>y�=zu����~&���i99���5�$�}���ۊ���v}:Ե7s3$Բ�s��8�����K�I}��F�3��V��E&�g�{|�����ϏG�;�ҍ���X�t��qv���sf�Yg.j�cS�u���{�)s�n)�1y���ξyN������;Ƀ���Y��|��z��u����˝n$?�����N�o.�|s�#'��s��$��^���	�I��S�-���,���|�o�=�,������z�kJ���`�&٘1��7r��ֹ�r�T2.���6�f97&��4�B�q(C�3�\��H�tٸ��لх �K��	�5IF�1�����6�Ĺ�f��d̚K�.`Y��jZ�l�B���+���%'>�׿�9��Nro���I�N�5�=����ӽ����V��>ۛ��?Fb��y4�d���7�g{kM)K��5��Y���G�2k���:�Z�����fy�n$��Hܜ3Fo�~γ�s�����������J�����땛GZbd6,�f��3i��5\�+��	��������ϿĒNr8��;�S��;U�{�%;���ľ�q��q�j}Ѽω�Ř���������LL'}_�}�w)���e���"�:rϳ������|�X�wZ[���#o����+�M�{���r{�u�kvW�k����yx^�#cY����K�\�ָ��6�yߧU��,���|e{zﻹoS7��f�y��\ۙ��mM͕�Wry����q�m��������������c0�A�� �a0�1�A� �ac0�A�� �a0�1�A�x��c0�A��5�z�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1����3�?���������<��<��<��<򪪪����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<��<��<��<��?��Ȉ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������c�1�������ǻ;���_nv�Bu�I&cѳv�Ù����͵7=4��9���,��)9�WXyOd�D������`ϊ�)p)p�%u5U6 ��g_����}y�dzh���qz��U{�Ȥ�f�����M}���O^�1zyrS�꧴s�{����ǯ��vN>�옒zC�i�N�ۜ��?v��z9�w��N�޹ֿn0Z|��s5۾?�'���Rm=��T�Ho��d2y�*8��x{-��Ggr�7kv���sS�q��S�S����"��K����$��&����P�+�EVӮOތ��}��?#Ͽ?xs��REt������Z{K���Os]���ّ:�������E�9�~3��f���?���Ց{wM�y��i�����%o��5�����I'9	'9<����k��N`�5-gn1��5���&�E�L��r�^K!��G���0�3�39Z�����\�0�hl&l&�AbL�ß�z맭bR��f&46���Ý콭-�ǝ����%���㧢�/SKZo_8u���a�Nsw/��'�1��!�~�yOI}w�<��ϓ�ω!�%���i�C��Lk�x�ȼ��;���yy�>I!������ۉ�ػ�+Qw�����������N��]'	����|���ɲ��>�p6�]M�nu�n�F�нw�rI9�Y$������n�������xx��&\��h��/�[k�?	���s?Lj��I9�5=�ϻػ��yNg�}��3�eosu���^Λ��<�q}�Oy�!��'�Z���T�]i-�i�jnT���$kÕ�GZbd6,�f��6���:4��{^�����=��`�ts�o�9|d�~U���}�r}��&99�w}���&$�'{�=�RH����#޷RoI����s����?��{�ǰ=�s�/��\��to�}������޿�W��W�$�y�]�wҿ��K�J���1��5؍�r
��qn�ָ��\�OϜ� G��ҝ���^��	S���5���1H�Ĭ�Z�w�3�4�ok����$�77���}�c��q������k����k��r��&1�׳�A99Ɏ�����k���G�Ӈo��;�7�<������ -�RWSUSb�um�j߃��~$�{Umy������q�nD7�f4L�j5������.}�+G5\=�ޒ��y��ͳW�P�'l��SɛZsU�mM�O�]���zRY�Q�6�_j5zz���$����trNr_>�4��f:$�4I��s��K��]ls��aHd]u�����Rr�nm�Z��ٰP������L����K�Z��i�3`�Z�0s�s��JQ�.#13��A�CD\�n᫱46n��ML�150]w������������w��y����̉�^K���[��Ru���}�T�y�ݯr{��1��g����/2G�L|��}����<��S'���#VM)���-�ק?I}�ي&��X���z�'���7��J7hf�%��M��v��Bj�1�ы,;�D��xII�'�'�1$��19�L��q�zz�?{�_��~���q� 9�Üi�m�<f��܍q�)qGƍ-�?24�^��������&�����>W�58���k�L������՟jN>&�b�ߚ��(گ���n���:��i4�Q=zG��RtD������{�zBgR�1�D�m���Z�v�+k|�W�|��xw��N�ǖ(������㜜�e�n��2}�&����94�����w\���9���a�1�0��B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B�������������u9��O���-?�=����Ś�|��&�����k��E�Q#������2zG�η�>v�f�֒�lض�]�6�����y���}��x��C�M��csk�G�ܛ϶=���I浖����[����{�Z|kz�r�I��}�q�Y�n���<|��w��������8���x�ə����5�6����������a�����4�b6-�Y���F�M����cz��E's8���9ć�5㚚\z�w/s5�.�6��SmϷ�!�.ǜ�kQuqwy�{�o}u<�4vM���y1���m�"j�>��}�|���r��7��d[�}��f�[F��E�tk2$��k$}�����������1�A� �ac0�A�� �a0�1�A� �ac0�A�� �fCSO��$ �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a3���������g����<��<��<��<�ʪ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<��<��<��<���0��K�;�����;�]>I<�9�0s��|���v��� �۝����%�s����nv�։'{��n�v��%���N�9�`s����O�O9�s��s�%�$ݷ9��;v�}�/zIc��s۷9פ�H�9���w��u�1�u��s���KZ֖9�݁���$���7m�w8�s��Z뮓�s��n��k�N�9�݀�ۜKKפ��s���s�׮�$�s��9��>KRI�ns{�v����^���9���ns�I$��s����I.�c��v��9뮖��,s��{��IkkZnۜ�p=��5ֵ�]'��/0.ݹ��Z$��s��۷8���I;�����;�]>I<�9�0s��|���v��� �۝����%�s��n��^�I#�g9ޒ]�H�9����s�]-kZX�;v�s���ִݷ9��{9�k�k��O9�^`]�s���I;��;v�nsM,�U+��GI�nV�¸��PĦ�cB�<2���sC��p��uo��fL�Mhc�b��R.�`c���,A�^&	�K��JVl�q3��FkDp8�mD���"�%������:� ����ݼ��ߋ9O�����}y���>w�t?o:�@��o?{�d�~�|t�j-?�R7�^�O���ɕ����=`�|���R7��#]����\ˉD��w�y�A�""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""#��9��������C��m�n65\���ƿ�Ei�����Y�.�]Zjg31��㩺��(�w��/���vO���Ց��#�%y��/v���b��^3����5����?y�߭�<mݤ�����>��<�u��ȳ1�ܖ7ݤ{�Z�m9��N����5���ǝ�mn�����<�W�v@���s�[���K�M-�лan!5n��h�J��u~���m���3�k����_���~�~���JO^mk��"�훙�sRE}7럴�_|�I�O�vG��0���N����|~$��F�53S������i����s}x��￞פ��[tA��l1�֗H1 ��=�z$���Oa���5$U�I�#�׸��ڳ��gz��.=}�1�j;�Uv������;LȌ|Ϣrw��j�\�����N�I��i����ӟ��I�9�r0� {���[I��ts����e9���߻Vy�<�	���6�i��Y�u��6-��a��樮^�Ood��q:�xuS�R@��^n�c��o��s/�[�?t�;_�s�'��"M�����vO=n#:#����SI����V~���Nď��Ş]f>:	$��/�g��$��u��z�~�������~����)���f���Nr}�Jx��1�ɸ�+�&1���1(j�:)3!��Z�W4 ����6]oX̆9�E�4scb��Qtk dËj׉�L.���JW`6#����R��p]f0��i��l[r
�n\[��7\���xJ7�	�1���m��[ε��I<��N���\q�sO�NE�o�-���Bk|�j���4Ϟ�Z�{"Oi�&L����Ϸ${��)$���|��B�~������l�
�:�ײ��ݝ_�珅�S�=�|�\	\�]����nʦ�9�X�y�Х�;^�߽1��vou�����=O�Ó6��/�Z�Ǐ�7ދc�a�q���7G���ٯ�7G]�����1���o��sI�W�ߋ�$���)��}g��޾�z�:7��կW���S�0�������y�����X�n�C�ּ;�ey��{��u���Svd�Ǥ<��Z��gr8��so�3>�]����s;���J�i�ie�=�I=%�'gY�������9��g�"H�	���v�^���|��GG'�w�Hs�?��vk"F��m#�M><��߅��{毯(/r��	I|��u[��Е�Ɩ������i�������ć����w��.e��}b�������&�}��N�G��Zh�ǥ���[�ɑoK�|��9ؖ�����o����t���{�����s���O�}�:&�w�=�I9��Nr_��3�UO�?�?����~k���S���o����{ �nA��l�nu��AB\��xw�>���wc���'��%�����;�u�:T����xɯw�}pi���g��zW�g����9���R{yӞ�|�}ߺ��}�b_�����l~�fI��:�ե�q��SKo	�\�ĒNI�p��������g	r�h�����tRfL*�ml
�kJē4��ւ�-e,��t]3a� lʲ�ٍ`LL�2aq��n\�$	�h�WB��q�0W#�j�0�f� h�P�r�7]uŝB�a.55��e6��^���������Ώ�#1��|�ݳ�ON���5y�|�����6�|~���SM������:��O��I9�����>��׽�ܷ���z�<g�v�V���"*�l�������oj�ȧqqk�5܃��]%Ź�[ �7&j~��9E����ݿ3}����k����Ns뻻�����G����'ĉ���\C_*�s"Ȟs'"��]8�%q���9:$��vwbq���z����S�N��c��M�/��L5�u��;/������S?����ߨ�D�f���E�/,�m�Tأ˜����>,ko��xY�F��Y���>�����T�w='�D��3�vWu�'�_���'[ȵ��k��%������������a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �� �� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac?���������������<��<��<��<��<��*�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<��<��<��:r!E�11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�0�Ō11cLX�jS���x�ꗓs���]η����q����6kL$�Q!��m7�̒+ɮ$�Ւr�ۃ]���N���O8�����k�M.��l�밲�j?��Ɏ_ߧ�cm����k�G���b{������U�w>��ly���dQ���!��_t�~k'Qwm�.�:�����}7��|1i餾�m�������w�8���u������_=�^��߼���.��n4�7]��isv73��e�_'�yR��NΏ��o~W�8��î�:����ב���k��q�\Y���$���qr��wkOo6{[o���},�$��3s�Ѿεu!2a��;��oqM�y��jE�c�	�zw\}�����Np����$��&���?��\8ӚK
�	r��p�.9���4.�́AqX����Z��(���A��:�4����f5	�0���1�h.���벅q�j�&v h�R��jك��-��]����R� ���{�]t�ۮzN$��ȜN8}�e��'G;9��c�(w��Os�<��#�y\�k��ԯ\�NdM�׸wq	I9�i�$�D��C���v�w��3ۥ�N�$;��������4o���3�6�g�+5����,�}|k��z[^��s�Sޭ?Lnк�3l�Zkf��R뱴�-	KW���Ϸ���곯]���_gw���zi��x���y'9+7�4��Q��#R��o��b��[$���7�^��%�7�=�|:/�R�����n�;�~�oN��1{꧞�����2�Y����E������=���x��1l�Y��r��t��l4���m�������`O{~���ӈ�x����釭{��q_s{�54c̓��dV�ٍ8��̯{�c_/�Z�Ǔ<��"�s�g2������Rq�y�>i��h�٤���߻����Y����9����l�k���2��2�e�F��������=��4�71�Ek�݈ps�&�=�ٙlǎ9�G�1=I�N�W���ncE�Lv� _a+�Ǧ��㯇��D�	'>Q�HM:���a5�a�-?��iiΎ�c����:9?O7R[�%�i���V�:]e��%�a��r���ȝ�G�S�'9N$�|�����嶢��[f�4�*�_r}=����]z�-ߗ��{������ݽ|ɷ��!�I��s�QL���o���*�9����ִ���]fCisNr�4l�%��:?ǜ�������pܼM%�3��XV��,a��2E��l�U�+�nL��]v�)Fd32�����XjQ�n�n�j��d��d:e���8@бt.Q�벅vaSV96�)��t�-�ܵ��.%cpiu��o4��^3332(�G��X��o��^�qq�%�z�j��z�<�}�D����I'9{��xf�I}�kZ�����ۯ�2�}k|����5��;>��Smɑ��z�7�q&񭗆ƺ��Vw7w�d��Ϻ�����y�>o;��P�� �Erֺ;T�β��C�.S��ڼql�M�o��~}$���0Ç^��K�_/�G仕��w�n.q�YMWs��9;����M�i�|L�<����s�}o=��~n,w�g�$�ֵ�޲������������i�ƃ4.���d�����R뱴�vI�E1��Ϻ���������N�GF��)���orj�ͤ���e�,kzFk��Y^>-�{���$�%���޻�v~�+�HP:߾�n�_u�H��ϗ�����9��3=�%Z���I_H���/5_�u�y���\ē��_+�5�Pu�t�˹qp�q�8kfu�y{�LO	;��~d��xxq������h��������|}��g���u�M�bf���rrĹ��KM�lb�'�JF��kMV���.��V�b_}��~q����e���|cy캜u�����QѲ��Yn�k�fWc�!��=�󟾿�z��w����O��z�y���Q���ǖI'9�Ä�ma���*�e�^��H�=͵�wz�>�,w�o��Z�����[��fg1�>ެ��s=&�����뿙�~p�(�Djj\XM=C!3��ۿ����_���� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�$ �ac0�A����6�a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A��/迢���?�������<��<��<��<��<�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<��<��<��<��?���G8�_�_�;��9�;��k]i�I'{��<�{���I%��M�s����s�׮���'��;��wp.ݹ�Ii$�v��n�39�Iiu�I��9�09��;Z�OzI;��9����zI/^�nۜ�n��ۜ�t��I<�9����;�I)$c���g9���M�i,s�n�v��w^�I$�9�3�s��I!$�s��{9�ֺ�ֵ���9���v�9%��M�s�� ��9%��]'{��<��s��k�=�$�s��ss��$�zI�ns���ns���w]$��{����$���s��=��;�I6����u�۷9�z�$�X�8���s�$��1�w8��;Z�KZ֞s����ۜ䖒I7m�v�3�䖗]t��s����s��������s�`=��w����&��v�ݹ���I�t��s��`�s����F9�^`�s��$�֒�9��n��u뤒Ic��0ow9���H�9�����k�-kZy�s���ns�ZI$ݷ9۰�s�Z[}���M!��5Ѩ\G,M��dt�&�+���77u���b�S,GB�8�`iF��eٍps d�.�cY�� �4\͇;)M�`j�7́���I]I`Zk���4t��m�]]�t)N����u��<k��$�7��I$��d}\�G�"�ߧ�0��|�3M˨���y;4��{�q�I�~nξ;�u���#������w��[7�f����k8ɭ.�|ȟ�9�����:��{��g��>�ϵ����kt��q+����P��uԱ�:���z��t8V3���w��3���+r{��73=>K�=���OM;����t�6�<^��c�k�g9�O5��]�w}�(��?I�=������r+�z�c�v����~#=9�sߺ֬
i(�����U��S����|�A��w�ֽ�$`��B4Q�1��m�Gg6�RZ�w G�{���_+��Ol���ߞ�9��Yv}�rGZV���Y��^�btr}.�������M���rn��I'�&�_|�Ƈ�f�%�k�s2rG��ĺ�~o{�~϶Ƹ׼��2%��)���O�|2|N�y�^y�7�$�OΧ����w���ݛ���//����������������>!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�F}��=����MzI�r&�����w{���z[���ƚ����J�}Y�h�hn$z��iQL��������4���{�S�{ca�1�0�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�B!�D"�BI��M&�iM�����D�̙(���g[�η����y�'���b�9��3)��b�pp�.���ߜ�����ۏ��|�'P�c�*w����Λ�To>��[����M�I'T�7�}���7q�Y������ǝ�~;ۿ|�N��s:��-����k2E�Og;�G���]{ژ{b�y�'9;띿����M!�u�u#P�qq2�hm�7&֖We3i7.�&�����A�q���Ҵ�S.�k�LD�CM6�IN��qsp9ٔՖ�sq�a��%.�\����fev6l�,�m��r�$�����|����~N��ܚs��;���ŏ�5q{��w�S�߈�O	�}uJ�s��ͯ$�����y���8|?�����t�g'�[���e�IYֱ!�����T��>k{'٫�I�����������znn��%�\�c7[����G�\���(�z�������G�:��o��^z��YΠ�����.��w���k��m��X���}z�)'���^C�'���\��zw���=��r~�~���?K����1>�L��A�$����Ժ�k;�i+}ʹݭ҆%ĬnK���B�s;Y������x~��׬����rk������S���J�'�kiZ�F��_X���>/����߬�$�'���/:��;�&��❝i�ۻM���֟'s$�zI6w���ϯ4�V�7��Z��{�X�S�ʈۘ�j��hY�@�k�߿w�\���L>�_χԦNI8
�7\'�o&q�w���S�$��s��F��O�;3�xisܼ�iLU�u�k���槽>�I}�i/�]�7���?M����Mi����旵����5��$��g�~��ƃ4.�;L�Z]�Z�v1�Y���r{�}�ׇ~�w�{��W:������G����8gZ���nv)'rM��y�޹<����Z�2,�sK;����r�>NI��f�V�fw/������w���?ĒNr{I'9<�O먼Ig4��[h�s��rY��mMrm[���f&��4	�Y�7R��WXA�q1uR��v�ɘ�a&dL��j�]�R�g-ʹٛ�f
�]	�d�1Ò��[�k0�݈iX�L�n����w՞���߽~��o��~M<�''=�wN^Ų��q�07���5ԓq��w7ˬ]};���%nfkDˬ9��m�Ǭ;[ڕ��]�f/_o_��s��=�^��s�����(�w�J�te,k�fV��Ś���l��3�������Z��{��v��_v$��i{���hֻ>�7�f&jo�f�9��q��u�j��7��_�u����g��#�f'���xnon��u?1F�5���yٷ�;zK�k��|�浙��I3Y��ߦ�����q�M�f�������������z��9��(�5�ٽs����������?O��DA� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� �a0�1�A� �ac0�A�� ��{{w����0/�)�?0)����F�6���E��h�Z-������������,h�cF�4XѢƌ�^=Q����cX�k�b�h�Z-�E�Q��ccb��ō���V�lV�ض�Ŵ��X�Z-�E��h�lX�ر��h�Z1���#d[Q�#j6Tm���6���-�E6M�d�6�O�6E�ڍ�ڋQTm���6�شZ-�E��h��h8����ϟ��y�y�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUW�I}�����8���I��o�5��FwY�<䛊�9��M;z��Ӕp��
\B��a�Z�/4��j<�ǧ5 nn��w�U�4g��MHmf;����n[����H^�~�]��~����7$��$ޗ|:ֽ���K��fN�i�r���i�.�����x<�H��۲�6�9��TvsB��h[$[��LL�5��4]�d��95��w��d��x��)�1��Vk-y۬ۼ�"��s=�u�_\�r�}�yI��Y���%�	�1�c�)��z��������=�>w��I'9	'9?u�*"�'�M�B�e.�ë5]�l�ɑ�Ck�c�M���.!�q��c�]`9���5v[�l�M�r�4���fo!�vj��&�5�Ĥ΅��!�%�IW���uߟ��<���hN�G���ch�WT�������N�ۮ~p�fG^k������q{��3��ˍ�kJ��s�~�Iɛû������HβI̘���e�|<�N��7�^�(��My��J�,2\B&�i�?�����߼�o����B2N���wש/�Gjɘ?uk&�kji�^��3���oےK�5���7d8vo�����ͧS$�w,���y�X���y2;�]e�2�5�3+pLb�V6�����5�c��}����Y&I�w�+����{�ky���9���ɴ��.�n�����3>��M�{�]W�\�g���$�7>�}��߿^�<?`�S��bKu��vn��L�h����c]\����.߻�ދ��fbȣ�=�L�Ľ1���I�޹o����nuw���}��&'������}��0a���DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr"#����DG""9Ȉ�DDr&�I����$�S�cgtws�.i�sϓ�?�R!K���a�Z�/4��%��?`���N�z���Q|S��7z�����_����z�Og���֝�������D�����of��K鿫5��Ed~���	)�������/����:�+ZW��&	�l���R霩�5�a��pd]Uf��Y�Mɤ,)G���J�+�5�1�H�u2�Sfl�hn%�̀k5��P��WSR�ic1.a��3&����4�;*#nc��;9��nF����՞}��n���[Ԛ��e�sYs5�{��rv^{�jE��+�l̞����`��gn�]_q�5�aٲ�$�F�������HxxN������/GPy�m��T�bm��Pn���f�]u6gg�gϟ����=tJ���<��=�����I�BI�G�m��޻��.H��dǼ��]�~^5g�h%�y3�3\����g����z�E4�y�y�� �}�����b�|�טPnĺi�e�K�8�� mSپ.w��=�=���m��;s������#|ߺ;��n�����I9���sR@���vؒK�^#�mf���d�(�3%�{w�gJ���+��k5��y�,�6»fd�Jb�aEq���v���^7������������F��'�"��9�~�_{���s�Ʋ���U���ڛ�I}�-<�$��V���M����{�D�뙃]u��f�ѵ�n�ƱJ6��>߱���:����do�����/�6cO�i��8��ou��9�>�}y��٫g�KI}��?{��Nݭ����#{#�Ѯo�>]����K�^[\U]]UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUW����DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��DD""��DB"!��O��s��$����N坣�����s��u��$���/0��;�I{�M�s���n��u��H��n�w�������䖏y$�w9�3g9�-.뤻��y���s��u��$���/0��;�I{�M�s���n��u��H��n�=��}�'�#�/09��;�I6���9�0ݹ���IK���ۜ�I!$��ns{�^�s��������9��{9�rKI$���8�g9�-.��s����9��Z{�Iy�r��ns�$��$ݷ9�݁v��w^�N뤏9�v���wޒ|�1�r���s���kZLs�� �ۜ�t�$��q�ݹ���I�v�7���;Z�KkZy�s�����$��I��s��fs����N�9�y���s��u��$���/0��;�I{�M�s���n��u��H��n�=��}�'�#�/09��;�I6���9�0ݹ���IK���ۜ�I!$��ns{�^�s��������9��{9�rKI$���8�\�:i��nY�D��2M��8�q����3�Pȩ���r�^K!�jQ�.���
s<31s�.)i��\�0�;	�	�F���:���蜱��f&46�&f��7�R%B����n����;�:�%��7�o�֝x��%ӣ��w��n#\�s�<w[�cx�/{g����8���^ffC�ߜ�׽�T;���Q�/}n}��>~��~�|#���Q��8f�ó��[7�F����=��s�\���Ǯ7��_|�sm;�ίE#܉��~3���r�MD�_|�dW�~���-���������_�y��鈃�d����<�OsM�I�}�DcA�-�&ҥ�m��Ꜷ,�´l�?��	�����{�k|��|��������}��s�
���u������$������������U�K)�:7��u��q�Mo��ܜ�/�k�9��{�ǯo|�w?uk�Pm��l���B��]j��޾=���|����ޛOq�����s��ܹ:�q�2Ǿ�U��4���=�.rk#ɞ�-������5ٱ%��Ѽ�;ǘ�rh�g�Ѭ��[�w<��[��ڶ»�a�c����=������_��'��j�k�����j��E��;9�>I$��ՒI�N��~��;Y�E��C~��u����>~f����{��@O����%B�z�s���կ�sI�h8��&���3�RU6�v�d��CsR�!q�x��\�jb�+���\�,a���L�8�`�&�9�Ĥ#�m���A�f��MG5�5�Zk�j�]�pV�\Q�3j|����[���,�N��Q7&�s���=�Wk|����m��.[��Ji$��*�57q���v�;O2��\}y�ݣ���[���3Z�8�F��o�_�B��"J��)�]��-�K.�V��e|�~��~���_��Ձ�[m���d����u�o_��<����:޸���뾿o�r��̎8�C\�&��j]�k���=�t���b��=Db���v��ݖ9�6��Պٸ2���:F���|��]{�\7�4�u�ƺsr�d���y�oڍ�9���%���\깳{[7tzdRN㗞]�wJn=�͛չ2Fk���񫮷�uߟ���!���K]t�i��n��eŬ3j�/�Z{�b�&�̓O~~�Z��t�x^4禖[�޺k@\Z���"�$��έ��۬�k��I/�[I}��׾�����}�n���sG}�����P�@�.�@�Ժm,4���9��jL����|O������{��ڵ?�=o�ϯ@�ԟ�&�222FN8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�p�qÎ8q�8��8�(�;?4ߌ�w��m��/��I�*wW�5���͸��,�5��6�5�}�b�����q�{���{�a��@�f�®q��r�u�Ά&�E�ZInn^'/�eթ����3�:LV�)2&�re.ekXC&���j�D��h:S5�ĥ��39�!ty�r\Xˠ]s*]�k���c��0ٶ`�d������=߾�μ�;��Ԓb޹���y޹9ɯ\qk..�]��Owy{:�NE$�B9�U�-�I�k�'r,���ۯ=�f{M��>m�����08�Ktѫ�+]�fu��Z�{뇣�k5��}��T�5��ߩ/�^��}m�I/�^��{�ܙ��zg5x�k=�^w=�9>��޶�F�Q�nI'�ɳ�پI���$��y��5�F�g$)�]�虩n�˰����soCh�!kr?y7�f8�9+��˛Z�Y�����o�����{�׍,�ҋj�.�B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!B�!u%�˝����͡�y���t��j�&��X��F�1e���|����u�9!���*'��`�Vm\;C*ق�lߵew�_���ڿ�*�w:�賛�T�_|���ط}��cȳ^��ɝn]woK����w&���5��|��_|��4�s$��Çcs�˧ێś��vd!�����]6�h��-�.����Ư^�����߳�t�Wy�sSx��{�s�I%�˾��Ǿ����z<�B/P�~�s���z��>B�W�xֳ_�齚�0�$�ț���j{z7��~m��z��$����'9>zS���VM�ܭs��6��%Y�E&xe5�������˭�����0�kC؛R��X�&X8�V�M`�t��T�f�lG���5��ຶ(l5�ۥ�f�it%b��6Vm��2�o�����zA��Oŉ�r��Mf���ܵ��=2ݬ�3�mc̛�7�{{�{m�5�s���1�c��s5��.�iH�{1G�$�֣���;��X�z���߰.�<�tY���C9�t+�c]t�r��ϖL�_�������gz��#���?���9��Vok�ᗼ��O�Ǯ�k]z�x�7��n�qe���w�&�{��z}i<o��>���9�<�O�};�e0Zl���]n�v��-�3�զ�~6Yp�{���Y^M$���6���������?���}��[�����O�S�F��ɶ�����y�MA�=Y�=�{��>O~/�ׅ�Oߕ}�*���IL�ёrl]٭��=�5��k�iL�a�+���-�nt�}����+��6�W~&>Dk���s��כY&I��4i��<�4�5�_=���mė�#�;���"}�S�"��μ�g�<�;J��M�6�6�U�ʮ�����F�}��~߯[����k8�sQ�z��o����G0��tާN<of�d�2L�oz��{�r��Σ��ks'{�ɳ9t�m�"K�}�M�hf&+ɸ��s��6��%��h:)3&r]��sJ�ē4����0Z�Y�aNh:.��ʐ6�eT��F�&&H0���n\��h.�Юk�kL�]ls�kR��j����7��K]t�i��n��cs43��y�^��ߋ７X�('�7�o�mh��7�柔�GW-���6Ws\zܑ���O5�^i���>y�K#ɺo���{��;��t������f��a%���iu#nk6���2{}#~���I}��t����杻���_���$�s��'9?���ܟ��T�.�m�Ù�]�Q�tָ�'�,QH��<�����ŭy��=śx�o��׽�z�d]�qm��u��K�:�t���c�4k���]R���ߺ����{�~����g����7�{�����vkn>�U+�;��'9<N�w^�s�F�y���oի�֞��޵s�bzU�oXo�ѥL~}�h�;]q5��7MCk���tsY�s����}5=���Vn��t��'2>��f��3oyx��dCz��1�)l{P\�5ʫo9���Ȧ�_����ye7�I}�Лפ�4���B�.��57�_���Y~���iL�cJW%��䱋lL��=��߻��k��x�Ÿ���]3b�.���57�᛼6�<�K��L��;��-�X�}�5�����W�NM�և���]��Gs�{ٚ������q5U�m˗��oo{ȿ�������"*�������������������=5
��%'`^}�])<d�^}�P��W�RS�
��R�h��*��$񪔽�A�O���ׯ����{��ϖ�c�|����Q����~��=��=�}��y���?�O���S��ÒD���������%��(���	G���n|�����-�}����?���χ���������}?7����v~��U������O�~�������*��E_��@���>/���C�������������@E[���ٟw�~�������_O}���OYއ>�O�u�����G�ƾ�u��ݻ�������s�}}�׻�U�>��׾_��<zu��?���������=�9XSS
i�Ņ1aM,)��1aL��
a&ҫ
j�
e
b�
e&�L)��)�<p�	0��0�R���0��aMB�C
i҆�SH��J����)�XSG吸S�SD����N¦�,)�SR��,)�SR�Җʌ)�S
`�)��)��S(����SXS)0���5XS+
iaM,)��4��,)��5XSS
baMS)�
haMSF�
haMS�aLF�0�V�aL�)��2\���z�ow˽��<zw���^c�������*��5pV��*�?���ߗ����y����~k�G�o���>����{|��z��E_�������~����O����@��}������z���~{�w����^���m�����~��~����6������������~�o���}�U����i���<~ϯϟ/�����U��P������~���>�������������<_ "�O��������W���F���m�ϡ�����c�z_���xOS�s{{���"�����'�y�/on~�=='�>���_�y{ýs��_��o��`W���)�/�����^8�w�g����:�5����o��o���~���O��s�w���?����I�U����Y��	��}��W�����=ߏ��������޷��=�7�g���^<���w�{������~_+���/����׏�}���*��x�۾/�_g�s�s���������^t��z�����<G��������}�hW�[��?Y��������������"����E_d��Ͽ������>��ݞ��﹟��>X�%��ן��ܑN$RA�@