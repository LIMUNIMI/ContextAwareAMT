BZh91AY&SYW��] ߀Py���������`
>��=��;ҥ.O�}�[5- ���Bz�A'��T�6�F&�d@0L@�F�	5�(      T��ꨏ�OP �      ?T�Ma4�a4�LF �M1 �D���ʃ�4ze i��ѣCF���)� ��Ld��� �!�=OS�e,@?@*�!h*ށ���I$!:o�Hp�8� �@9��N�H\��E���4QN�%RD���|�R-��@>TG"">�b�G�3�WH�,r���5�K8xHԣD��aW9�w�ܩ)g�r�t�z������ۅ��'0'0YdD
�",��@H
�"
�"
�/x���4��D�H�4f�����<`R//����~��Z��)c=��n�M0,���SR��h�����#��6�H�xy�-N�km���\� švrWg$�  '1\�����)J�*R�k\�rC�ar�r*x7L�R1I�`���ہ[y�;������k���86,�KX�
Ta�
� �Z"�{��$ah�(�IU���b�	�2�y[8���$�����lkz�uƷL�V*��I^ 	��( ��Se^Q[���F%y�aŧ�il�{[G�s�^F���j�J'�
s�	���+7|\CZ]�u�I$�#HIQ:P�:��µ�3߮�$a��S��z7y�k�F3ۋgJ�TU�)\�*�uɥs��c �NM���I$�I���TN�'N� 3��D���m���%-�$Ix��4fg|�sma�����4}L)�\��V�nr,�02.y��9x��M'qlE�$�I$�LeL�%	ҌVy�����BF���V�rSr�� Hk�+FU�<`[vV�/J���N���         �<� ���z=ؤŔ�)_M�CαL�{Y���%�K�|��%�9�c��P��BEIU.]i��ԛ5$�+U~�05����݀)��\*|V�S8�&�Eфmz�HH�ZO����D�Q3��`�ܵ.@r���kPED�"� $�� �<If}�ci��'�� �z&�;��Bp�	" �A֔��L=���oY}�76@s� �B
|���t�*/��ˏ��XC7�uZ'rJ��� ��U^=z"�ȒT�y�� ��UI�1��ݻ��i� y��_�u	��R�ڈt"kAL�#�^A	
�ƒE6�k���ê�ީ�*��������I�wD�@)rb.5)�:�H�%��.�C�Q8��W�v5J
�P���JS���6 �(R���L`<�#���֖���chP��q����IP���H�j� �v D��Yr�� "  
�K�@ D @*��1'�VUW(�.���e
�J~wLx9�*..��]m R�U�P$#�)J�s	�xqܬ���.p2Wx�h�	�l�n]V��$큀�X>i�]���'�<�ݿ��(EJ��y�G��_Kw�C�>�Y�Ow@(��*/m���{���S�*�v�l�'�6%;�O�5�y��;W�HL���b}�_-����H%{��S�"�q@o�:��|މ=�9���_0��R�`yW`
Y6�P�D�
"y+�D�Ԧ�H�,
�!],!T����+��t<�"��Bd%���@ �*)�0��Ѕ���(�T�R�?�2P�/V��f@)=�4<��9�W�
iJw���4�8"`��gd��z�4`fCP�����ɜ�7���uF�Ū�=�������*���">�#}'֯P ���\.j|��	�5�tC����r�����0�_��D�59�(�s,w�x.��5��հ���ܾ�aj�)2�N� S)6��]�[F���hG�v��>�SJ[r�9�T�^��*�k���vm�D�VkZ�TL�U�
d縻��^���P�
qEM���Q~W/��,�	r��hYj�QS4�:����)����