BZh91AY&SY\��l ^߀Py���������`]�v��IU��  � �`�2��JhDI��4F��� � 9�#� �&���0F&jH��h�I��4�    h9�#� �&���0F&
� �&Ɓ��)<MM��� hh�4�4�HG�m	%��dI��c�Q���Z��h�f��q�Tĩ%R�]),���T���JTO���B^�:�U�4�yt#�n�&X#��a//e�[�]}�	�3bj2��n��ߎ�:��vme<<�E7��ے0���C!���5 �`1��'}Z�=�|lc1�T���F�7��]f�Bl��~�x������������Fԏ��5���Fs��b���&�fa��<��1�&<�ZNA��{��͊� �1C4�"�၄��D�ޮ�e�uX�20%�d����&B XX�ĴLW��6dGkGv�Y+����J)���ÉQg#��1�c�Q!�ɡ�q�a��[j.ڞbw�M'\�2������u,�J"*c�4�C���ɚ�+�I5w��q�9�:���.��ΉrF��sn��4�|4皙|\)�g%�h�A�[����#����I)�����|`�+9�
7���AYu��,�oD�?(*pSقK��>4���*/\J�I	�M��a���=���֎pk����eNH'w/��3�s��)���.��&K�i�q�;�ATԨ�TJ(��⓷!���iPD�X�h�R��#,@�ɡ�E���2��Fl�\�j�󦀙w�#&Rv0����b�(c�C<C ��ߔ���ȅ�f�B�ƃ4<�S'ȡ�.�o��3���3�o���Fi� <����;��!QQ��b"g28a����LxK2)��}��-����XKQ�|tgI�UUUUd�ו�����9�z���O2>�I�Iꓲl�~1i%)c�Ng�[�>��������*�B��\�v�]ߤ��خ�ܙᾧ�t�)J0E�agA�IbV_*F�L�������k~Y��Q���8e�o�opT��H�-��!�C�>��t�JiX#L��#K��E�״%ܢ�Ցb�09�gFt�r��v5���d�'��郙(�JR�U�K]��ٚ)ǜ��bz��N�IEvVΓ���90�������8�=�S�%%"�	a��s�H�b��G?��c�03N��6��
W��������ùS�6*�uI���wNF��{�rtԊV��}:J<͋���jԟ��˟�K�}"0v���=�J�Q�W�~��ʗ�⹌�}�̗71�k^�&��;$5T���}X�faag�%F݌)Q$��
�?�2x�3^ɒ]Y���j��R?���a2�)&�P1��N�Ij���3�-�
hVM$�R��ʞ-$+��GBzOkg����{W��'�f<>�����$�<c��+����uv诰�z��Լ�w����t�� �I�|�όU%RU%T�N���}%���k�����F�yc&��*��EG/B�+�Vlu\��Gt�����f�l50��ZN�YlL�� �j5�L�)�Q��
U��A�i
�9�g�E'-Ƨ6�Q������1�f�^����c�IR~��y��$խd�К�͟;�7/%���]v?<q�'I�T3���R�-}!�t�!����"�(H.O̶ 